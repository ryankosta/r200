`ifndef _mux_vh_
`define _mux_vh_
`include "mux2w32.v"
`include "mux4w32.v"
`include "mux8w32.v"

`endif
