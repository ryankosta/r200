`ifndef _alu_vh_
`define _alu_vh_ 
`include "not32.v"
`include "or32.v"
`include "xor32.v"
`include "and32.v"
`include "and32s.v"
`include "adder32.v"
`include "shifter/mshifter32.v"
`include "shifter/shifter32b1.v"
`include "shifter/shifter32b2.v"
`include "shifter/shifter32b4.v"
`include "shifter/shifter32b8.v"
`include "shifter/shifter32b16.v"
`include "mux.vh"

`endif
