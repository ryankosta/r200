`ifndef _shifter_vh_
`define _shifter_vh_
`include "mshifter32.v"
`include "shifter32b1.v"
`include "shifter32b2.v"
`include "shifter32b4.v"
`include "shifter32b8.v"
`include "shifter32b16.v"

`endif
