`ifndef _comp_vh
`define _comp_vh
//comparitors
`include "comp1b.v"
`include "comp4b.v"
`include "comp16b.v"
`include "comp32bs.v"
//conditional logic
`include "condsel.v"
`include "condgen.v"

`endif
