module r200wb(
	wbsel,
	dmem_out,
	alu_res,
	pcp4,
	reg_win //instrn [11:7]
);
//input
input wire [1:0] wbsel;
input wire [31:0] dmem_out;
input wire [31:0] alu_res;
input wire [31:0] pcp4;
//output
output wire [31:0] reg_win;


mux4w32 wbselector( //select which data written into register
	.a(alu_res),
	.b(dmem_out),
	.c(pcp4),
	.d(32'b0),
	.sel(wbsel),
	.out(reg_win)
);

endmodule
