`ifndef _mux_vh_
`define _mux_vh_
//5 bit
`include "alu/mux2w5.v"
//32 bit
`include "alu/mux2w32.v"
`include "alu/mux4w32.v"
`include "alu/mux8w32.v"

`endif
