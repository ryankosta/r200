`ifndef _comp_vh
`define _comp_vh

//comparitors
`include "comp/comp1b.v"
`include "comp/comp4b.v"
`include "comp/comp16b.v"
`include "comp/comp32bs.v"

//conditional logic
`include "comp/condsel.v"
`include "comp/condgen.v"

`endif
